----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    05:43:08 12/30/2016 
-- Design Name: 
-- Module Name:    ANDP - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ANDP is
    Port ( zeroIn : in  STD_LOGIC;
           branchIN : in  STD_LOGIC;
           andOut : out  STD_LOGIC
			  );
end ANDP;

architecture Behavioral of ANDP is

begin
	andOut<= zeroIn and branchIN;

end Behavioral;

