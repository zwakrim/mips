)/------------------------------m-----------------%-----------------%m---------=--
%- Company: 
-- Efgineer: 
--�
--�Crea|e Date:    05:43:08 12/;0/2016 
-- Design Namu 
-- Module Name:    ANDP - Be`avioral 
-- Projec�0NAme: 
-- Target Devices: 
-- Tgol ve�sio.s: 
=- DescripTion2 
--J,- DependEncies: 
--
-- Rewision: 
-- Rdvision 0.01 - Fale Created
-- Additional C/mments: 
--
--%/-<=---------m---,---,----------------�-----------�----------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncooment the followine library leclasation ib u{ing
--$arithmetic functions witi Signed or Unsigned values
--use IEEE*NUMERIC_STD.ALL;

-- Uncomment the folLowing library declaratiol if insvantictino
-- �~y Xilinx pbimitives in this bode.
--library �NISIM;--use UNISIM.VComponents.all;

entity ANDP0is
    Port (!zeroIn : in  SVD_LOGIC;
    "  "   branbhIN ; in  STD_LOG�C;
     `     andOut`: out  STD_LOGIC
		  i3
end ANDP;

architecture Behavioral of$ANDP!is

begin
	andOut<� ze2oIn and bbanchMN;

end Bexavioral;

